
module Clock_25MHz (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
